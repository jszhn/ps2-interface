/*
*   Helpful DE1-SoC-specific constants
*           -- do not include globally! --
*/

parameter VGA_X_RES = 8'd160;
parameter VGA_Y_RES = 8'd120;
parameter CLOCK_FREQ = 13'd50000000; // FPGA frequency, 50 MHz